2�d d        d   * ��  Cxor2�   �����   �����   �����   ���� XOR     ��  Cpin�   �����   ����0 0                  ��   �����   ����1 1                   ��   �����   ����1 1                  �_  �����  l���l  �����  ���� XOR     �_  ����r  ����1 1                  �_  x���r  x���1 1                   ��  ~����  ~���0 0                  ��  Cswitch%   ����U   ����"   ����B   ���� X0     �%   ����3   ����1 ��                 �%   ����3   ����0 ��                  �U   ����G   ����0 1 X0"   ����        �!   $���Q   ���   E���?   3��� Y0     �!   $���/   $���1                    �!   ���/   ���0                     �Q   ���C   ���0 0 Y0   E���        �!   ����Q   ����   ����A   ���� Cin     �!   ����/   ����1                    �!   ����/   ����0                     �Q   ����C   ����1 1 Cin   ����        ��  Cand2�   ����   �����   -����   ��� AND     ��   ����   ���0 0                  ��   ����   ���1 1                   ��   	����   	���0 0                  ��   �����   �����   �����   ���� AND     ��   �����   ����1 1                  ��   �����   ����1 1                   ��   �����   ����1 1                  ��   ~����   Z����   �����   ~��� AND     ��   r����   r���0 0                  ��   f����   f���1 1                   ��   l����   l���0 0                  ��  Cor3  ����F  ����  ����4  ���� OR     �  ����  ����0 0                  �  ����  ����1 1                  �  ����  ����0 0                   �E  ����7  ����1 1                  �  Z���  *���  C���;  1��� X1    �  *���  8���1                    �  *���  8���0                     �  Z���  L���0 0 X1  h���        �P  X���\  (���f  A����  /��� Y1    �P  (���P  6���1                    �\  (���\  6���0 Z                   �V  X���V  J���1 1 Y1O  f���        �<  Y���H  )���R  B���r  0��� X2    �<  )���<  7���1 0                  �H  )���H  7���0                     �B  Y���B  K���1 1 X2;  g���        �u  ^����  .����  G����  5��� Y2    �u  .���u  <���1                    ��  .����  <���0                     �{  ^���{  P���0 1 Y2t  l���        ��  `����  0����  I����  7��� X3    ��  0����  >���1                    ��  0����  >���0                     ��  `����  R���0 0 X3�  n���        ��  e����  5����  N���  <��� Y3    ��  5����  C���1                    ��  5����  C���0                     ��  e����  W���0 1 Y3�  s���        ��  ����3  �����  ����)  ���� XOR     ��  ����  ����1 1                  ��  ����  ����0 0                   �2  ����$  ����1 1                  ��  >���2  ����  P���'  >��� AND     ��  2����  2���1 1                  ��  &����  &���0 0                   �1  ,���#  ,���0 0                  ��  ����5  �����  ����*  ���� AND     ��  �����  ����1 1                  ��  �����  ����0 0                   �4  ����&  ����0 0                  ��  ����7  ����   ����,  ���� AND     ��  ����  ����0 0                  ��  ����  ����0 0                   �6  ����(  ����0 0                  �l  E����  !���y  W����  E��� AND     �l  9���z  9���1 1                  �l  -���z  -���1 1                   ��  3����  3���1 1                  �m  ����  ����z  ����  ��� AND     �m  ����{  ����1 1                  �m  ����{  ����0 0                   ��  �����  ����0 0                  �o  �����  ����|  �����  ���� AND     �o  ����}  ����1 1                  �o  ����}  ����0 0                   ��  �����  ����0 0                  �  @���E  ���  R���:  @��� AND     �  4���  4���1 1                  �  (���  (���0 0                   �D  .���6  .���0 0                  �  ���E  ����  ���:  ��� AND     �  ����  ����1 1                  �  ����  ����1 1                   �D  ����6  ����1 1                  �  ����H  ����  ����=  ���� AND     �  ����  ����0 0                  �  ����  ����1 1                   �G  ����9  ����0 0                  %�v  �����  �����  �����  ���� OR     �v  �����  ����0 0                  �v  �����  ����0 0                  �v  �����  ����0 0                   ��  �����  ����0 0                  %��  ���  �����  ���  ��� OR     ��  �����  ����1 1                  ��  �����  ����0 0                  ��  �����  ����0 0                   �  ����  ����1 1                  %�}  ����  �����  ����  ��� OR     �}  �����  ����0 0                  �}  �����  ����1 1                  �}  �����  ����0 0                   ��  �����  ����1 1                  ��  Cprobe�  �����  �����  �����  ����  S0     ��  �����  ����0 0 S0�  ����          z��  �����  �����  �����  ����  S1     ��  �����  ����1 1 S1�  ����          z�  ����  ����  ����5  ����  S2     �  ����  ����0 0 S2
  ����          z��  �����  �����  �����  ����  S3     ��  �����  ����0 0 S3�  ����          �m  |����  X���z  �����  |��� XOR     �m  p����  p���1 1                  �m  d����  d���0 0                   ��  j����  j���1 1                  �`  �����  ����m  �����  ���� XOR     �`  ����s  ����0 0                  �`  ����s  ����1 1                   ��  �����  ����1 1                  ��  }���  Y����  ����	  }��� XOR     ��  q����  q���1 1                  ��  e����  e���1 1                   �  k���  k���0 0                  ��  ����=  ����  ����3  ���� XOR     ��  ����  ����1 1                  ��  ����  ����0 0                   �<  ����.  ����1 1                  �s  �����  ^����  �����  ���� XOR     �s  v����  v���1 1                  �s  j����  j���1 1                   ��  p����  p���0 0                  z��  ����  ����                        ��  �����  ����1 1                    ��   �����   ����                       ��   �����   ����0 0                  ��   �����   ����1 1                   ��   �����   ����1 1                  ��  d����  @����  v����  d��� XOR     ��  X����  X���1 1                  ��  L����  L���1 1                   ��  R����  R���0 0                  ��  j���7  F���   |���-  j��� XOR     ��  ^���  ^���0 0                  ��  R���  R���1 1                   �6  X���(  X���1 1                  �^  o����  K���k  �����  o��� XOR     �^  c���q  c���0 0                  �^  W���q  W���1 1                   ��  ]����  ]���1 1                  - ��  Cnet0  ��  Csegment�   �����   �������   �����   ������j   �����   ������U   ����j   ������j   ����j   �����j   r���j   ������   ���j   ������   ����   ������   r���j   r������   r����   r�����U   ����U   ����   "   ��0       ��1  ��_  ����_  �������   ����_  �������   �����   ������_  ����_  ����    ��1  ��_  x���_  x�����_  x���_  �������   ����_  ������Q   �����   ������Q   ����Q   ������Q   f���Q   �������   ����Q   �������  �����   �������   �����   �������   �����   �������   �����   ������Q   f����   f�����Q   ����Q   f������   f����   f�����Q   ����Q   ������Q   �����   �������   �����   �������   �����   �������  �����  �������  �����  L������  L����  L������  ����Q  �������  R����  R�����U  ����Q  ������Q  ����Q  W�����^  W���Q  W�����^  W���^  W������  �����  R��� 	 � #  � � �   ��0  ��  	����   	������   	����   	�����  ����  ������  ����  	��� '   ��Z       ��1  ��  ����  �������   �����   �������   ����  ���� (    ��0  ���   ����  ������  ����  �������   l����   l������   l����   ���� )  $ ��Z       ��Z       ��1  ��E  ����E  ������E  �����  �������  �����  �������  �����  �������  �����  �������  �����  �������  �����  -������  -����  -������  2����  -������  2����  2������  -����  �������  �����  �������  �����  �������  �����  ���� D H L  * ��Z       ��0  ��  Z���  Z�����  ���  Z�����  Z���  Z�����  �����  �������  �����  �������  �����  ������  ����  �����  ����  ������  &����  ������  &����  &�����  ���  �����  ����  ������  �����  ������  �����  ���� E I Q  . ��1  ��V  X���V  X�����V  X����  X������  X����  X��� �  2 ��1  ��n  p���n  ������2  ����n  ������2  ����2  ������n  p���m  p�����m  p���m  p��� �  F ��0  ��v  ����v  ,�����1  ,���v  ,�����1  ,���1  ,�����v  ����v  ���� l  J ��0  ��4  ����v  ������4  ����4  ������v  ����v  ���� m  N ��0  ��v  ����v  ������6  ����v  ������6  ����6  ������v  ����v  ���� n  R ��0  ���  �����  �������  �����  �������  �����  �������  ����o  ������o  ����o  ������o  ����o  �������  �����  ������`  �����  �������  �����  �������  ����m  ������m  ����m  ������m  ����m  ������`  ����`  �������  �����  ���� ] Y  o ��Z       ��0  ���  ~����  ~������  �����  �������  ~����  ~������  �����  ~��� |  
 ��1  ��  ����-  ������-  ����-  ������  ����  ������-  ����  ������  ����  ������  ����  ������-  ����-  �������  ����-  ������-  ����  ������-  ����-  ������  ����  �������  �����  �������  �����  �������  �����  ���� i e �  t ��0  ���  p����  p������  �����  p������  �����  �������  p����  p������  p����  p������  �����  ���� �  � ��1  ���  j����  j������  �����  �������  �����  j��� ~  � ��Z       ��0  /��  k���  k�����
  ����m  ������  ����  k�����  k���  k�����  ����  ���� �  � ��1  ��B  Y����  Y������  �����  Y�����B  Y���B  Y������  ����`  �������  �����  ������`  ����`  �������  C����  �������  ����o  ������o  ����o  ������o  ����o  �������  �����  C������  C���l  C�����l  9���l  C�����l  9���l  9��� � \ T  6 ��0  ��{  ^���{  ^�����{  ^����  ^������  ^����  ^��� �  : ��1  ���  q����  ����0���  �����  �������  q����  q��� �  � ��1  ���  �����  3������  3����  3������  3����  3������  �����  ���� q  V ��0  ���  �����  �������  �����  �������  �����  �������  �����  ���� r  Z ��0  ���  �����  �������  �����  �������  �����  �������  �����  ���� s  ^ ��0  ���  `���K  `�����K  ����K  `������  `����  `�����K  �����  �������  �����  �������  �����  ������K  )���K  ������K  ����  ������  ����  ������  ����  ������K  ����K  )�����K  )���  )�����  (���  )�����  (���  (��� � h a  > ��0  ���  e����  e������  e���(  e�����(  e���(  c�����^  c���(  c�����^  c���^  c��� �  B ��1  ��s  v���s  ������<  ����s  ������<  ����<  ������s  v���s  v��� �  � ��0  ��}  ����}  .�����D  .���}  .�����D  .���D  .�����}  ����}  ���� v  b ��1  ��}  ����}  ������D  ����}  ������D  ����D  ������}  ����}  ���� w  f ��0  ��}  ����}  ������G  ����}  ������G  ����G  ������}  ����}  ���� x  j ��1  ���  �����  �������  �����  �������  �����  �������  �����  ���� �  y ��1  ��s  j���s  j�����r  j���s  j�����r  j���r  >�����r  >���  >�����r  >���r  ������r  ����r  ������r  ����  ������  ����  ������  ����  ������  4���  >�����  4���  4������  ]����  ]������  �����  ]������  ]����  ]������  ����(  ������(  ����r  ���� � d `  � ��1  ���  e����  e������  e���
  e�����
  ,���
  e�����
  ����
  ,�����
  ,���l  ,�����l  -���l  ,�����l  -���l  -���T��
  ����
  �������  ����
  ������m  ����m  ������6  X���G  X�����G  ����G  X�����6  X���6  X�����G  �����  ���� � U X  � ��0  ���  �����  �������  �����  ������7  �����  ������7  e���7  ������7  ����7  ������7  ����7  �������  ����7  �������  �����  �������  �����  �������  �����  ������7  e���n  e�����n  d���n  e�����n  d���m  d�����m  d���m  d������  R����  R������  �����  R������  R����  R������  ����7  ���� M P �  � ��0       ��1  ���   �����   �������   �����   �������   �����   �������   �����   �������   /����   �������   �����   �������   /���^   /�����^   ����^   /�����^   �����   ������^   ����^   ������   ���^   ������   ����   �����^   ����^   �����^   �����   ����     � ��0 
 ��Q   ���U   �����U   c���U   �����Q   ���Q   �����U   c���
   c�����
   ����
   c�����
   ����p   ������p   ����p   ������p   �����   �������   �����   �������   �����   ���� �     17702