2�d d         �   ��  Cinput_signal:   ����p   y���G   ����`   ���� A       ��  Cpinp   ����b   ����1 1 AG   ����         ��  Csignal    0 ��   0 ��  0 �X  0 �   0 ��  0 ��  0 �x  0 �@  1 �  1 ��  1 ��  1 �`	  1 �(
  1 ��
  1 ��  1 �9   ���o   ���F   )���_   ��� B       �o   ���a   ���1 1 Bo   ���         �    0 ��   0 ��  0 �X  0 �   1 ��  1 ��  1 �x  1 �@  0 �  0 ��  0 ��  0 �`	  1 �(
  1 ��
  1 ��  1 �6   ����l   ����C   ����]   ���� C       �l   ����^   ����1 1 Cl   ����         �    0 ��   0 ��  1 �X  1 �   0 ��  0 ��  1 �x  1 �@  0 �  0 ��  1 ��  1 �`	  0 �(
  0 ��
  1 ��  1 �:   9���p   '���G   K���a   9��� D       �p   0���b   0���1 1 Dp   >���         �    0 ��   1 ��  0 �X  1 �   0 ��  1 ��  0 �x  1 �@  0 �  1 ��  0 ��  1 �`	  0 �(
  1 ��
  0 ��  1 �� 	 Cinverter�   ����  p����   ����
  ���� NOT     ��   �����   ����1 1                   �  ����   ����0 0                  L��   ����  �����   ����  ���� NOT     ��   �����   ����1 1                   �  ����  ����0 0                  ��  Cand2�  ����  �����  ,����  ��� AND     ��  ����  ���1 1                  ��  ����  ���1 1                   ��  ����  ���1 1                  S��  ����:  j���  ����/  ���� AND     ��  ����  ����0 0                  ��  v���  v���1 1                   �9  |���+  |���0 0                  S��  ����B  ����  ����7  ���� AND     ��  ����  ����1 1                  ��  ����  ����0 0                   �A  ����3  ����0 0                  S�Y  i����  E���f  {����  i��� AND     �Y  ]���g  ]���0 0                  �Y  Q���g  Q���1 1                   ��  W����  W���0 0                  S��  ���C  ����  ���8  ��� AND     ��  ����  ����0 0                  ��  ����  ����1 1                   �B  ����4  ����0 0                  ��  Cor2�  H����  $����  Z����  H��� OR     ��  <����  <���0 0                  ��  0����  0���0 0                   ��  6����  6���0 0                  h�(  ����l  ����5  ����Z  ���� OR     �(  ����;  ����0 0                  �(  ����;  ����0 0                   �k  ����]  ����0 0                  ��  Cprobe�  �����  �����  ����  ����  F     ��  �����  ����0 0 F�  ����           ��  Cnet1  ��  Csegment�  �����  ����v��   �����   ����v�l   ����l   ����v��   �����   ����v�l   �����   ����v��   �����   Q���v�Y  Q����   Q���v�Y  Q���Y  Q��� Q b  ) t�Z       t�1  v�r  ����  ���v�o   ���o   ���v��  ����  ���v�o   ���r  ���v�r  ����r  ���v��  �����  ����v��  ����r  ���� U ]   t�1  v��  �����  0���v�p   0����  0���v�p   0���p   0���v��  ����  ���v��  �����  ����v��  ����  ����v��  �����  ���� V f  ; t�1  v�p   ����p   ����v��   �����   ����v�p   �����   ���� N   t�Z       t�1  v��  v����  ���v��  ����  ���v��  ����  ���v��  v����  v��� Z  W t�0  v�  ����  ����v��  �����  ����v�  �����  ����v�  ]���Y  ]���v�  ����  ]���v�Y  ]���Y  ]��� Y a  O t�0  v�  �����  ����v�  ����  ����v��  �����  ���� ^  R t�0  v��  �����  W���v��  W����  W���v��  W����  W���v��  �����  ���� e  c t�0  v��  <����  |���v�9  |����  |���v�9  |���9  |���v��  <����  <��� j  [ t�0  v��  0����  ����v�B  �����  ����v�B  ����B  ����v��  0����  0��� k  g t�0  v�(  ����(  ����v�A  ����(  ����v�A  ����A  ����v�(  ����(  ���� o  _ t�0  v�(  ����(  6���v��  6���(  6���v��  6����  6���v�(  ����(  ���� n  l t�0  v��  �����  ����v�k  �����  ����v�k  ����k  ����v��  �����  ���� s  p   17702