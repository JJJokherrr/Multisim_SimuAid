2�d d           ��  Cclock'   !���]   ���4   3���U   !���
 Ck       ��  Cpin]   ���O   ���0 1 Ck4   3���        �� 
 CDflipflop�   �����   #���                       ��   I����   I���0 0                  ��   a����   a���1 1                  ��   �����   y���1 1                  ��   #����   1���1 1                   ��   a����   a���1 1                  ��   I����   I���0 0                  ��  ����A   ���                       ��  F���  F���0 0                  ��  ^���  ^���1 1                  �  ����  v���1 1                  �   ���  .���1 1                   �A  ^���3  ^���1 1                  �A  F���3  F���0 0                  �r  �����  "���                       �r  H����  H���0 0                  �r  `����  `���0 0                  ��  �����  x���1 1                  ��  "����  0���1 1                   ��  `����  `���1 1                  ��  H����  H���0 0                  ��  Cswitch�   �����   ����                       ��   �����   ����1 X                  ��   �����   ����0 Z                   ��   �����   ����1 0                  �~   �����   ����                       �~   �����   ����1                    �~   �����   ����0                     ��   �����   ����1 1                  ��  ����  ����                       ��  �����  ����1                    ��  �����  ����0                     �  ����  ����1 1                  ��  ����  ����                       ��  �����  ����1                    ��  �����  ����0                     �  ����  ����1 0                  �V  �����  ����                       �V  ����d  ����1                    �V  ����d  ����0                     ��  ����x  ����1 0                  �d  �����  ����                       �d  ����r  ����1                    �d  ����r  ����0                    ��  �����  ����1 1                  ��  Cprobe
  ����  f���  ����9  ����  Qc     �  f���  t���1 1 Qc  ����          4�j  ����~  `���w  �����  ����  Qb     �t  `���t  n���1 1 Qbw  ����          4��  �����  b����  ����
  ����  Qa     ��  b����  p���1 1 Qa�  ����          ��  Cor2�  o����  K���                       ��  c����  c���0 0                  ��  W����  W���1 1                   ��  ]����  ]���1 1                  ;�M   r����   N���                       �M   f���`   f���1 1                  �M   Z���`   Z���1 1                   ��   `����   `���1 1                  ��  Cand2P   �����   ����                       �P   ����^   ����1 1                  �P   ����^   ����1 1                   ��   �����   ����1 1                  D�M   Z����   6���                       �M   N���[   N���1 1                  �M   B���[   B���1 1                   ��   H����   H���1 1                  4�m   :����   ���z   L����   :���  Ck     �w   ���w   (���0 0 Ckp   ���           ��  Cnet1  ��  Csegment�   �����   ����Q��   �����   ����Q��   �����   ����Q��   �����   ���� 	   O�1  Q��   #����   ����Q��   �����   ����Q��   �����   ����Q��   #����   #��� 
  # O�1 
 Q�  f���  a���Q�  a���  a���Q��   a����   a���Q�  f���  f���Q��   a���  a���Q�  a���  ����Q�M   B���   B���Q�   ����   B���Q�M   B���M   B���Q�   ����  ���� 6 K   O�1  Q�  ����  ����Q�  ����  ����Q�  ����  ����Q�  ����  ����   ' O�1  Q�   ���  ����Q�  ����  ����Q�  ����  ����Q�   ���   ���   + O�1  Q�t  `���t  ^���Q�[  ^���t  ^���Q�A  ^���A  ^���Q�t  `���t  `���Q�A  ^���[  ^���Q�[  ^���[  ����Q�P   ����>   ����Q�>   ����>   ����Q�P   ����P   ����Q�>   ����[  ����Q�>   ����>   N���Q�M   N���>   N���Q�M   N���M   N��� 8 F J   O�1  Q��  �����  ����Q��  �����  ����Q��  �����  ����Q��  �����  ����   / O�1  Q��  �����  ����Q��  "����  "���Q��  "����  "���Q��  �����  "���   3 O�1  Q��  b����  `���Q��  `����  `���Q��  `����  `���Q��  b����  b���Q��  `����  `���Q��  `����  ����Q�P   ����I   ����Q�I   ����I   ����Q�P   ����P   ����Q��  �����  ����Q�I   �����  ����Q��  �����  W���Q��  W����  W��� : G >   O�0  Q��   I����   ���Q�w   ����   ���Q�]   ���]   ���Q��   I����   I���Q��   ����  ���Q��  F����  ���Q��  F����  F���Q��  ���r  ���Q�r  H���r  ���Q�r  H���r  H���Q�]   ���w   ���Q�w   ���w   ���Q�w   ���w   ���    N   O�0  Q�A  F����  F���Q��  �����  F���Q�A  F���A  F���Q��  �����  ����Q��  c����  ����Q��  c����  c��� =   O�1  Q��   a����   `���Q��   `����   `���Q��   `����   `���Q��   a����   a���   C O�1  Q��   ����4  ����Q�4  ����4  ����Q��   �����   ����Q�4  ����M   ����Q�M   f���M   ����Q�M   f���M   f��� A  H O�1  Q��   H����   H���Q��   !����   H���Q��   H����   H���Q��   !���   !���Q�   U���   !���Q�   U���M   U���Q�M   Z���M   U���Q�M   Z���M   Z��� B  L O�1  Q��  ^����  ]���Q��  ]����  ]���Q��  ]����  ]���Q��  ^����  ^���   ? O�0  Q��   I����   I���Q��   �����   I���Q��   I����   I���Q��   ����A  ����Q�A  b���A  ����Q�A  b���r  b���Q�r  `���r  b���Q�r  `���r  `���      17702