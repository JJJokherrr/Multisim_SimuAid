5�d d           ��  Cclock  ����7  w���                         ��  Cpin7  ����)  ����0 1                  �� 
 CDflipflop�  8���  ����                       ��  �����  ����0 0                  ��  ����  ���1 1                  ��  8����  *���1 1                  ��  �����  ����1 1                   �  ����  ���0 0                  �  �����  ����1 1                  ��  9����  ����                       ��  �����  ����0 0                  ��  ����  ���0 0                  ��  9����  +���1 1                  ��  �����  ����1 1                   ��  ����  ���1 1                  ��  �����  ����0 0                  �x  ;����  ����                       �x  �����  ����0 0                  �x  ����  ���0 0                  ��  ;����  -���1 1                  ��  �����  ����1 1                   ��  ����  ���1 1                  ��  �����  ����0 0                  ��  Cswitch�  W����  K����  i����  W��� ClrN    ��  K����  K���1 Z                  ��  W����  W���0 Z                   ��  Q����  Q���1 1 ClrN�  _���        ��  �����  �����  �����  ���� PreN    ��  �����  ����1 ��                 ��  �����  ����0                     ��  �����  ����1 1 PreN�  ����        ��  Cprobe!  ����5  ����.  ����P  ����  Qc     �+  ����+  ����0 0 Qc$  ����          $��  ����  ����  ����'  ����  Qb     �  ����  ����1 1 Qb�  ����          $��  �����  �����  ����  ����  Qa     ��  �����  ����1 1 Qa�  ����          ��  Cor2M  $����   ���                       �M  ���`  ���0 0                  �M  ���`  ���0 0                   ��  ����  ���0 0                  ��  Cand3�  ,����  ���                       ��  &����  &���0 0                  ��  ����  ���0 0                  ��  ����  ���1 1                   ��  ����  ���0 0                  +�V  "����  ����                       �V  ���i  ���0 0                  �V  
���i  
���1 1                   ��  ����  ���1 1                  ��  Cand2U  (����  ���                       �U  ���c  ���0 0                  �U  ���c  ���0 0                   ��  ����  ���0 0                  :��  ���  ����                       ��  �����  ����0 0                  ��  �����  ����1 1                   �  �����  ����0 0                  $��  �����  �����  �����  ����  CLK     ��  �����  ����0 0 CLK�  ����           ��  Cnet1 
 ��  Csegment�  8����  Q���G��  Q����  Q���G��  Q����  Q���G��  8����  8���G��  Q����  Q���G��  Q����  9���G��  9����  9���G��  Q����  Q���G��  ;����  Q���G��  ;����  ;��� 	     E�1 
 G��  �����  ����G��  �����  ����G��  �����  ����G��  �����  ����G��  �����  ����G��  �����  ����G��  �����  ����G��  �����  ����G��  �����  ����G��  �����  ���� 
    # E�0  G��  ����D  ����G�D  ���D  ����G��  �����  ����G�x  ���x  ���G�x  ���D  ���G��  �����  ����G��  X����  ����G��  ����  ���G��  X����  ���G��  ����  ���G��  X����  X���G��  X���2  X���G�2  ����2  X���G�2  ����U  ����G�U  ���U  ����G�U  ���U  ���  3 =   E�1  G��  ���  ���G�  ����  ���G��  ����  ���G�  ����  ���� (   E�0  G�  ���+  ���G�+  ����+  ���G�  ���  ���G�+  ����+  ����G�+  ����+  ����G�  ���  ���G�  ���  N���G�U  ���D  ���G�D  N���D  ���G�U  ���U  ���G��  N���  N���G�D  N����  N���G��  N����  ����G��  �����  ����G��  �����  ���� & < @   E�0  G��  ����  ���G��  ����  ���G��  ����  ���G��  ����  ���   / E�0  G�x  ����x  ����G��  ����x  ����G�x  ����x  ����G��  �����  ����G��  �����  ����G��  �����  ����G��  �����  ����G��  �����  ����G��  �����  ����G�7  �����  ����G��  �����  ����G��  �����  ����G�7  ����7  ����G�7  ����7  ����    D   E�0  G��  �����  ����G��  7����  ����G��  �����  ����G��  7����  7���G��  &����  7���G��  &����  &��� 2   E�1  G�  ����  ���G��  ���  ���G��  ����  ���G�  ����  ���� 4   E�0  G��  ����  ���G��  �����  ���G��  ����  ���G��  ����M  ����G�M  ���M  ����G�M  ���M  ��� .  5 E�1  G��  ���7  ���G�7  v���7  ���G��  ����  ���G��  v���V  v���G�V  
���V  v���G�V  
���V  
���G�7  v����  v���G��  v����  ����G��  �����  ����G��  �����  ����G��  �����  ����G��  �����  ����G��  ����  ���G��  ����  ����G��  �����  ���� 8 A *   E�0  G�  ����&  ����G�&  ����&  ����G�  ����  ����G�&  ����<  ����G�<  ����<  ���G�M  ���<  ���G�M  ���M  ��� -  B E�0  G��  ����  ���G��  �����  ���G��  ����  ���G��  �����   ����G��   ����   ����G��   ���V  ���G�V  ���V  ��� 7  > E�1  G��  ����  ���G��  ����  ���G��  ����  ���G��  ����  ���   9   17702