2�d d            ��  Cinput_signal&   ����\   ����3   ����L   ���� A       ��  Cpin\   ����N   ����1 1 A\   ����         ��  Csignal    0 �d   0 ��   0 �,  0 ��  1 ��  1 �X  1 ��  1 �&   ]���\   K���3   o���L   ]��� B       �\   T���N   T���1 1 B\   b���         �    0 �d   0 ��   1 �,  1 ��  0 ��  0 �X  1 ��  1 �"   ����X   ����/   ����I   ���� C       �X   ����J   ����1 1 C/   ����         �    0 �d   1 ��   0 �,  1 ��  0 ��  1 �X  0 ��  1 ��  Cand2  ����V  ����  ����K  ���� AND     �  ����   ����1 1                  �  ����   ����1 1                   �U  ����G  ����1 1                  "�  `���R  <���  r���G  `��� AND     �  T���  T���1 1                  �  H���  H���1 1                   �Q  N���C  N���1 1                  ��  Cand3  ����O  ����  ���A  ���� And     �  ����  ����1 1                  �  ����  ����1 1                  �  ����  ����1 1                   �N  ����@  ����1 1                  ��  Cor2  ]���K  9���  o���9  ]��� OR     �  Q���  Q���1 1                  �  E���  E���1 1                   �J  K���<  K���1 1                  ��  Cxor2�  �����  |����  �����  ���� XOR     ��  �����  ����1 1                  ��  �����  ����1 1                   ��  �����  ����0 0                  6�  =���R  ���  O���H  =��� XOR     �  1���!  1���0 0                  �  %���!  %���1 1                   �Q  +���C  +���1 1                  "�  j���S  F���  |���H  j��� AND     �  ^���  ^���1 1                  �  R���  R���1 1                   �R  X���D  X���1 1                  ��  Cprobef  M���z  -���s  _����  M���  F2     �p  -���p  ;���1 1 F2i  -���          C�n  y����  Y���{  �����  y���  F2S     �x  Y���x  g���1 1 F2Sm  Y���           ��  Cnet1  ��  Csegment\   ����\   ����J�  ����  ����J�i   ����\   ����J�i   ����i   E���J�  E���i   E���J�  E���  E���J�i   ����i   ����J�  ����i   ����J�i   ����  ����J�i   ����i   ����J�  ����  ���� $ 4 -   H�Z       H�1  J�  ����  ����J�  �����   ����J��   T����   ����J��   T���\   T���J�  T����   T���J��   T����   ����J��   �����   ����J��   �����   ^���J�  ^����   ^���J�  ^���  ^���J�  T���  T���J�\   T���\   T���J�  �����   ����J�  ����  ����J�  ����  ���� % @ ( .   H�1  J�  H���  H���J��   H���  H���J��   ����  ����J�  ����  ����J�X   ����X   ����J��   Q���  Q���J�  Q���  Q���J��   �����   Q���J��   �����   H���J�X   ����X   ����J��   �����   ����J��   ����X   ���� ) / 3   H�1  J�Z  K���J  K���J�J  K���J  K���J�  R���  R���J�Z  R���  R���J�Z  R���Z  K��� A  5 H�1  J�U  ����g  ����J�g  ����g  ����J�U  ����U  ����J��  �����  ����J��  �����  ����J�g  �����  ���� 8  & H�1  J�Q  N���h  N���J�h  ����h  N���J�Q  N���Q  N���J�h  �����  ����J��  �����  ���� 9  * H�0  J��  �����  ����J��  1����  ����J��  �����  ����J�  1���  1���J�  1����  1��� <  : H�1  J�N  �����  ����J��  %����  ����J�N  ����N  ����J�  %���  %���J�  %����  %��� =  0 H�1  J�Q  +���Q  +���J�p  -���p  -���J�p  +���p  -���J�Q  +���p  +��� E  > H�1  J�x  X���z  X���J�R  X���R  X���J�R  X���x  X���J�x  X���x  Y���J�x  Y���x  Y��� G  B   17702