2�d d         d    ��  CMuxesA  b����  ����                       ��  CpinA  J���O  J���Z Z             0    �A  :���O  :���0 0             1    �A  *���O  *���0 0             2    �A  ���O  ���1 1             3    �A  
���O  
���0 0             4    �A  ����O  ����1 1             5    �A  ����O  ����1 1             6    �A  ����O  ����Z Z             7    �Y  ����Y  ����0 0             A0    �c  ����c  ����1 1             A1    �m  ����m  ����1 1             A2     ��  ����w  ����1 1             Z                 ��  CplusV�   �����   ����                          ��   �����   ����1 1                  ��  Cground�   k����   S���                          ��   k����   ]���0 0                  ��  Cswitch	  ����9  ����  ����7  ���� A0    �9  ����+  ����1                    �9  ����+  ����0                     �	  ����  ����0 0 A0�  ����        �	  ����9  w���  ����7  ���� A1    �9  w���+  w���1                    �9  ����+  ����0 0                   �	  }���  }���1 1 A1�  ����        �  L���5  @���  ^���3  L��� A2    �5  @���'  @���1                    �5  L���'  L���0                     �  F���  F���1 1 A2�  T���        ��  Cprobe�  *����  
���                        ��  
����  ���1 1                    ��  R���  ���                       ��  @����  @���1 1             0    ��  4����  4���0 0             1    ��  ����  $���0 0             A0     �  7���  7���1 1             Z                 ��  ����#  ����                       ��  �����  ����0 0             0    ��  �����  ����1 1             1    �  ����  ����0 0             A0     �#  ����  ����0 0             Z                 ��  H����  <����  Z����  H��� I0     ��  H����  H���1                    ��  <����  <���0                     ��  B����  B���1 0 I0�  P���        ��  �����  �����  �����  ���� I1     ��  �����  ����1                    ��  �����  ����0                     ��  �����  ����0 0 I1�  ����        #�  W���'  7���   i���A  W���  Y0     �  7���  E���1 1 Y0  7���          #�  ����.  ����'  ����H  ����  Y1     �$  ����$  ����0 0 Y1  ����          ��  -���  ����  ���V  ��� CROSS    ��  �����  ���1                    �  ����  ���0                     �  -���  ���0 0 CROSS�  ;���         ��  Cnet0 
 ��  Csegment�   *����   :���B�A  :����   :���B�A  :���A  :���B��   k����   k���B��   *���A  *���B��   
����   *���B�A  *���A  *���B��   
���A  
���B��   k����   
���B�A  
���A  
���      @�Z  B�A  J���2  J���B�2  Y���2  J���B�A  J���A  J���    @�Z  B�A  ����A  ����B�A  ����A  ����    @�1 
 B��   �����   ���B�A  ����   ���B�A  ���A  ���B��   �����   ����B��   ����A  ����B��   �����   ����B�A  ����A  ����B��   ����A  ����B��   ����   ����B�A  ����A  ����  
 	   @�0  B�Y  ����Y  ����B�	  ����Y  ����B�	  ����	  ����B�Y  ����Y  ����    @�1  B�c  ����c  }���B�	  }���c  }���B�	  }���	  }���B�c  ����c  ����    @�1  B�m  ����m  F���B�  F���m  F���B�  F���  F���B�m  ����m  ����   " @�1  B��  �����  ����B��  
����  ����B��  �����  ����B��  
����  
��� %   @�1  B�  7���  7���B�  7���  7���B�  7���  7��� 9  * @�0  B�$  ����#  ����B�$  ����$  ����B�#  ����#  ���� ;  / @�1  B��  @����  B���B�g  B����  B���B��  B����  B���B��  @����  @���B��  B���g  B���B�g  B���g  ����B��  ����g  ����B��  �����  ���� ' -  3 @�0  B��  �����  4���B��  4����  4���B��  4����  4���B��  �����  ����B��  �����  ����B��  �����  ����B��  �����  ���� ( ,  7 @�0 	 B�  -���r  -���B�r  ����r  -���B�  -���  -���B�r  ����  ���B��  ����  ���B��  ����  ���B�r  ����  ����B�r  ���r  ����B�  ����  ���� ) .  ?   17702