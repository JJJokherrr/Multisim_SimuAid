2�d d          ( ��  CclockN  Y����  G���[  k���~  Y��� CK       ��  Cpin�  P���v  P���0 1 CK�  ^���        �� 
 CDflipflopy  �����  0����  �����  ���� D     �y  V����  V���0 0 CKm  d���        �y  n����  n���0 0 D3i  |���        ��  �����  ����1 1 S�  ����        ��  0����  >���1 1 R�  0���         ��  n����  n���1 1 Q3�  |���        ��  V����  V���0 0 Q3'�  d���        �x  �����  2����  �����  ���� C     �x  X����  X���0 0 CKg  f���        �x  p����  p���0 0 D2h  ~���        ��  �����  ����1 1 S�  ����        ��  2����  @���1 1 R�  2���         ��  p����  p���0 0 Q2�  ~���        ��  X����  X���1 1 Q2'�  f���        �M  �����  3���Z  ����s  ���� B     �M  Y���[  Y���0 0 CK>  g���        �M  q���[  q���0 0 D1=  ���        �o  ����o  ����1 1 Sk  ����        �o  3���o  A���1 1 Rk  3���         ��  q����  q���0 0 Q1�  ���        ��  Y����  Y���1 1 Q1'�  g���        �*  ����n  0���7  ����P  ���� A     �*  V���8  V���0 0 CK  d���        �*  n���8  n���0 0 Q0'  |���        �L  ����L  ����1 1 SH  ����        �L  0���L  >���1 1 RH  0���         �n  n���`  n���1 1 Q0n  |���        �n  V���`  V���0 0 Q0'n  d���        ��  Cand4  ����`  ����                       �  ����*  ����1 1 Q3  ����        �  ����*  ����1 1 Q2'
  ����        �  ����*  ����1 1 Q1'
  ����        �  ����*  ����0 0 Q0'
  ����         �_  ����Q  ����0 0                  ��  Cand3  W���a  3���                       �  Q���+  Q���0 0 Q2  _���        �  E���+  E���0 0 Q1  S���        �  9���+  9���1 1 Q0  G���         �`  E���R  E���0 0                  ��  Cor2�  �����  ����                       ��  �����  ����0 0                  ��  �����  ����0 0                   ��  �����  ����0 0                  ��  Cand2�  �����  ����                       ��  �����  ����0 0 Q2�  ����        ��  �����  ����1 1 Q1'�  ����         ��  �����  ����0 0                  4��  ����  [���                       ��  s����  s���0 0 Q0'�  ����        ��  g����  g���0 0 Q2�  u���         ��  m����  m���0 0                  )��  ;����  ���                       ��  5����  5���1 1 Q2'�  C���        ��  )����  )���0 0 Q1�  7���        ��  ����  ���1 1 Q0�  +���         ��  )����  )���0 0                  ��  Cor3  ����\  ����                       �  ����+  ����0 0                  �  ����,  ����0 0                  �  ����+  ����0 0                   �[  ����M  ����0 0                  )�  ����G  ����                       �  ����  ����0 0 Q3'�  ����        �  ����  ����0 0 Q1�  ����        �  ����  ����0 0 Q0'�  ����         �F  ����8  ����0 0                  )�6  }���z  Y���                       �6  w���D  w���0 0 Q3'$  ����        �6  k���D  k���1 1 Q1'$  y���        �6  _���D  _���1 1 Q0&  m���         �y  k���k  k���0 0                  /�{  �����  ����                       �{  �����  ����0 0                  �{  �����  ����0 0                   ��  �����  ����0 0                  ��  CswitchW  �����  ����d  ����}  ���� S     �W  ����e  ����1                    �W  ����e  ����0                     ��  ����y  ����1 1 S�  ����        V�Q  ����  ���^  "���x  ��� R     �Q  ���_  ���1                    �Q  ���_  ���0                     ��  
���s  
���1 1 R�  ���        ��  Cprobe�  �����  n����  �����  ����  Q3     ��  n����  |���1 1 Q3�  n���          _��  �����  o����  �����  ����  Q2     ��  o����  }���0 0 Q2�  o���          _��  �����  p����  �����  ����  Q1     ��  p����  ~���0 0 Q1�  p���          _�d  ����x  n���q  �����  ����  Q0     �n  n���n  |���1 1 Q0f  n���          4�s   �����   ����                       �s   �����   ����0 0 Q3'a   ����        �s   �����   ����1 1 Q2'a   ����         ��   �����   ����0 0                  4�'  ����k  ����                       �'  ����5  ����0 0 Q2  ����        �'  ����5  ����1 1 Q0  ����         �j  ����\  ����0 0                  4�'  Z���k  6���                       �'  N���5  N���0 0 Q2  \���        �'  B���5  B���0 0 Q1  P���         �j  H���\  H���0 0                  4�,  ����p  ����                       �,  ����:  ����0 0 Q2  ����        �,  ����:  ����1 1 Q0  ����         �o  ����a  ����0 0                  4��  ����2  ����                       ��  �����  ����0 0 Q3'�  ����        ��  �����  ����1 1 Q2'�  ����         �1  ����#  ����0 0                  )�n   O����   +���                       �n   I���|   I���0 0 Q3'\   W���        �n   =���|   =���1 1 Q1'\   K���        �n   1���|   1���0 0 Q0'\   ?���         ��   =����   =���0 0                  )�w  �����  ~���                       �w  �����  ����1 1 Q3g  ����        �w  �����  ����1 1 Q2'e  ����        �w  �����  ����1 1 Q0g  ����         ��  �����  ����1 1                  )�+  ���o  ����                       �+  ���9  ���1 1 Q3  ���        �+  ���9  ���1 1 Q2'  ���        �+  ����9  ����0 0 Q0'  ���         �n  ���`  ���0 0                  /��   ����   ����                       ��   �����   ����0 0                  ��   �����   ����0 0                   �  ����  ����0 0                  B��  �����  w���                       ��  �����  ����0 0                  ��  �����  ����0 0                  ��  }����  }���0 0                   ��  �����  ����0 0                  B��  �����  ����                       ��  �����  ����0 0                  ��  �����  ����0 0                  ��  �����  ����1 1 Q3�  ����         ��  �����  ����1 1                  "�:  ����~  ����                       �:  ����H  ����0 0 Q3'(  ����        �:  ����H  ����0 0 Q2*  ����        �:  ����H  ����1 1 Q1'(  ����        �:  ����H  ����0 0 Q0'(  ����         �}  ����o  ����0 0                  _�  ����)  ����"  ����V  ����  R_NS     �  ����  ����0 0 R_NS  ����          _��  �����  �����  �����  ����  Y_NS     ��  �����  ����1 1 Y_NS�  ����          _��  �����  �����  ����  ����  G_NS     ��  �����  ����0 0 G_NS�  ����          _��  �����  �����  ����  ����  R_EW     ��  �����  ����1 1 R_EW�  ����          _�t  �����  �����  �����  ����  Y_EW     �~  ����~  ����0 0 Y_EWn  ����          _�'  ����;  ����4  ����m  ����  G_EW     �1  ����1  ����0 0 G_EW   ����          4�,  a���p  =���                       �,  U���:  U���0 0 Q2  c���        �,  I���:  I���0 0 Q1  W���         �o  O���a  O���0 0                  $ ��  Cnet0          ��1  ��  Csegment�  n����  n������  n����  n��� a $ � � �   ��1    	     Z ��1    
     ^ ��0    I N i y } �   ��0  ���  o����  p������  o����  o������  p����  p���	 c + 6 ; m q u � �   ��0  ���  p����  p������  p����  p������  q����  p������  q����  q��� e , ? J r �   ��0  ��_  ����_  �������  �����  �������  �����  ������_  �����  ���� 1  ( ��0  ���  E���`  E�����`  E���`  E������  �����  �������  �����  E��� 2  . ��0  ��  �����  �������  �����  ������  ����  ���� D  8 ��0  ���  m����  m������  �����  m������  m����  m������  ����  ������  ����  ������  ����  ���� E  < ��0  ��  ����  )������  )���  )������  )����  )�����  ����  ���� F  A ��0  ��F  ����F  ������{  ����{  ������{  ����F  ���� S  L ��1    % > j z � �   ��1    & 7 O ~ �   ��0     ' : K  � �  ! ��1       ��0  ��y  n���y  �������  ����y  �������  �����  ������y  n���y  n���   3 ��0  ��x  p���x  ������[  ����x  ������[  ����[  ������x  p���x  p���   G ��0  ���  �����  �������  4����  �������  �����  �������  4���M  4�����M  q���M  4�����M  q���M  q���   U ��1       ��0  ��{  k���{  j�����{  ����{  ������{  ����{  k�����{  k���y  k�����y  k���y  k��� T  Q ��0  ���   �����   �������   �����   �������   �����   ���� �  k ��0  ���   =����   =������   =����   =������   �����   �������   �����   =��� �  � ��1  ��n  n���n  n�����n  n���n  n��� g - @ P n v �    ��0  ��  ����  ������  ����  ������  ����  ���� �  � ��1  ���  �����  �������  �����  �������  �����  ���� �  � ��0  ���  �����  �������  �����  ���� �  � ��1  ���  �����  �������  �����  �������  �����  ���� �  � ��0  ��}  ����}  ������~  ����}  ������~  ����~  ������}  ����}  ���� �  � ��0  ��1  ����1  ������1  ����1  ������1  ����1  ���� �  { ��0  ���  �����  ������j  �����  ������j  ����j  �������  �����  ���� �  o ��0  ��j  H���{  H�����{  ����{  H�����j  H���j  H�����{  �����  �������  �����  ���� �  s ��0  ���  }����  �����n  ����  �����n  ���n  ������  }����  }��� �  � ��0  ���  �����  ������o  �����  ������o  ����o  �������  �����  ���� �  w ��0  ��o  O���~  O�����~  ����~  O�����o  O���o  O�����~  �����  �������  �����  �������  �����  ���� �  �   17702