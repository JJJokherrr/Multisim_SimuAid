2�d d         d    �� 
 CFullAdderR  x����  &���                       ��  Cpint  &���t  4���0 0                 ��  &����  4���1 1                 ��  F����  F���1 1                   �R  F���`  F���1 1                  �~  x���~  j���0 0                  ��  s���  !���                       ��  !����  /���0 0                 ��  !����  /���0 0                 �  A����  A���1 1                   ��  A����  A���0 0                  ��  s����  e���1 1                  ��  n���G  ���                       �  ���  *���1 1                 �%  ���%  *���0 0                 �G  <���9  <���0 0                   ��  <����  <���0 0                  �  n���  `���1 1                  �  i���i  ���                       �3  ���3  %���1 1                 �G  ���G  %���0 0                 �i  7���[  7���0 0                   �  7���  7���0 0                  �=  i���=  [���1 1                  ��  Cxor2�  ����  �����  ����  ���� XOR     ��  �����  ����1 1                  ��  �����  ����0 0                   �  ����  ����1 1                  �  ����K  ����  ����A  ���� XOR     �  ����  ����1 1                  �  ����  ����1 1                   �J  ����<  ����0 0                  �>  �����  ����K  ����x  ���� XOR     �>  ����Q  ����1 1                  �>  ����Q  ����1 1                   ��  ����s  ����0 0                  �Z  �����  ����g  �����  ���� XOR     �Z  ����m  ����1 1                  �Z  ����m  ����1 1                   ��  �����  ����0 0                  ��  Cswitch  c���  3���  q���.  _��� X3    �  3���  A���1 X                  �  3���  A���0                     �  c���  U���1 0 X3  q���        ,�S  e���_  5���i  N����  <��� Y3    �S  5���S  C���1                    �_  5���_  C���0                     �Y  e���Y  W���1 0 Y3R  s���        ,�  m���  =���!  V���A  D��� X2    �  =���  K���1                    �  =���  K���0                     �  m���  _���1 1 X2
  {���        ,�G  j���S  :���]  S���~  A��� Y2    �G  :���G  H���1                    �S  :���S  H���0 Z                   �M  j���M  \���1 0 Y2F  x���        ,��  o����  ?����  X���  F��� X1    ��  ?����  M���1                    ��  ?����  M���0                     ��  o����  a���0 0 X1�  }���        ,�'  i���3  9���=  R���^  @��� Y1    �'  9���'  G���1                    �3  9���3  G���0                     �-  i���-  [���1 1 Y1&  w���        ,��  p����  @����  Y����  G��� X0    ��  @����  N���1                    ��  @����  N���0                     ��  p����  b���0 1 X0�  ~���        ,��  n���  >���  W���/  E��� Y0    ��  >����  L���1                    �  >���  L���0                     ��  n����  `���0 0 Y0�  |���        ,��  ?����  3����  Q����  ?��� Cin    ��  3����  3���1 Z                  ��  ?����  ?���0 Z                   ��  9����  9���1 1 Cin�  G���        ��  Cprobe3  ����G  h���@  ����a  ����  S3     �=  h���=  v���1 1 S36  h���          Q�  ����%  n���  ����?  ����  S2     �  n���  |���1 1 S2  n���          Q��  �����  p����  �����  ����  S1     ��  p����  ~���1 1 S1�  p���          Q�t  �����  w����  �����  ����  S0     �~  w���~  ����0 0 S0w  w���          Q��  [����  ;����  m����  [���  Cout     ��  ;����  I���0 0 Cout�  ;���           ��  Cnet1  ��  Csegment  A���  F���^�R  F���  F���^�R  F���R  F���^�  A���  A���    \�0  ^�G  <���G  A���^��  A���G  A���^��  A����  A���^�G  <���G  <���    \�0  ^�i  7���i  <���^��  <���i  <���^��  <����  <���^�i  7���i  7���    \�0  ^��  �����  n���^��  n����  n���^��  n����  n���^��  �����  ����   L \�1  ^�,  ����0  ����^�  ����  ����^�  ����,  ����^�,  ����,  &���^��  &���,  &���^��  &����  &���    \�0  ^�t  &���t  p���^��  p���t  p���^��  p����  p���^�t  &���t  &���   H \�1  ^�Z  ����Z  ����^�Z  ����Z  ����^�9  ����Z  ����^��  �����  ����^��  �����  ����^��  �����  ����^��  9����  ����^��  9����  9���^��  9����  9���^��  9����  F���^��  F����  F���^��  F����  F���^��  ����  ����^�  ����  ����^�  ����  ����^�  ����  ����^�  ����9  ����^�9  ����9  ����^�>  ����9  ����^�>  ����>  ���� )   ! %  P \�0  ^��  !����  o���^��  o����  o���^��  o����  o���^��  !����  !��� 
  @ \�1  ^�  ����  i���^�-  i���  i���^�-  i���-  i���^�  ����  ���� "  D \�0  ^�J  ����J  ���^�J  ����J  ����^�J  ����  ���^��  !����  ���^��  !����  !���   # \�1  ^�>  ����>  j���^�M  j���>  j���^�M  j���M  j���^�>  ����>  ���� &  < \�0  ^��  �����  ���^��  �����  ����^��  ���%  ���^�%  ���%  ���^�%  ���%  ���   ' \�1  ^�  m���  ���^�  m���  m���^�  ���  ���   8 \�1  ^�Y  e���Y  ����^�Z  ����Y  ����^�Z  ����Z  ����^�Y  e���Y  e��� *  4 \�0  ^��  �����  ����^��  ����  ����^��  �����  ����^��  ���G  ���^�G  ���G  ���^�G  ���G  ���   + \�1  ^�3  ���3  c���^�  c���3  c���^�  c���  c���^�3  ���3  ���   0 \�1  ^�=  h���=  i���^�=  h���=  h���^�=  i���=  i��� S   \�1  ^�  n���  n���^�  n���  n��� U   \�1  ^��  p����  s���^��  p����  p���^��  s����  s��� W   \�0  ^�~  w���~  w���^�~  x���~  x���^�~  w���~  x��� Y   \�0  ^�  7���  ;���^��  ;���  ;���^��  ;����  ;���^�  7���  7��� [     17702