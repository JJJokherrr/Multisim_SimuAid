2�d d        d    �� 	 Cinverterw  ]����  9����  o����  ]��� NOT     ��  Cpinw  K����  K���0 0                   ��  K����  K���1 1 Yuxuan Zhang�  Y���        ��  Cswitch   W���K   K���K   _����   M��� Switch1     �   W���)   W���1 Z                  �   K���)   K���0 ��                  �K   Q���=   Q���0 0 Switch1K   _���        �   ����K   ����(   ����l   ���� Switch 2     �   ����)   ����1                    �   ����)   ����0                     �K   ����=   ����0 0 Switch 2K   ����        ��  Cand2�   ]���   9����   o����   ]��� AND     ��   Q����   Q���0 0                  ��   E����   E���0 0                   ��   K����   K���0 0                  ��  Cnand2�   ����  �����   �����   ���� NAND     ��   �����   ����0 0                  ��   �����   ����0 0                   �  �����   ����1 1                  ��   ����  ����                       ��   �����   ����0 0                  ��   �����   ����0 0                   �  �����   ����1 1                   ��  Cnet0 
 ��  Csegmentx   Q����   Q����K   Q���K   Q����K   Q���x   Q����x   Q���x   ������   ����x   ������   Q����   Q�����   �����   ������   �����   ������   �����   ������   �����   ����     
 �0 
 �K   ����K   ������   �����   �����K   �����   ������   �����   E�����   E����   E�����   E����   E�����   �����   ������   �����   ������   �����   ������   �����   ����      �0  �w  K���w  K����w  K����   K�����   K����   K���      17702