2�d d           ��  Cclock   1���L   ���                
         ��  CpinL   (���>   (���0 1                  �� 
 CDflipflop�   �����   ���                       ��   D����   D���0 0                  ��   \����   \���1 1                  ��   �����   t���1 1                  ��   ����   ,���1 1                   ��   \����   \���1 1                  ��   D����   D���0 0                  �  ����G  $���                       �  J���  J���0 0                  �  b���  b���0 0                  �%  ����%  z���1 1                  �%  $���%  2���1 1                   �G  b���9  b���1 1                  �G  J���9  J���0 0                  ��  Cswitchw   �����   ����                       �w   �����   ����1                    �w   �����   ����0                     ��   �����   ����1 1                  �w   ����    ���                       �w   ����   ���1                    �w    ����    ���0                    ��   ����   ���1 1                  ��  ����  ����                       ��  �����  ����1                    ��  �����  ����0                     �  ����  ����1 1                  ��  ���  ���                       ��  ����  ���1                    ��  ����  ���0                     �  ���  ���1 1                  �V  �����  ����                       �V  ����d  ����1                    �V  ����d  ����0                    ��  ����x  ����1 1                  �c  ����  ���                       �c  ���q  ���1                    �c  ���q  ���0 ��                  ��  ����  ���1 1                  ��  Cprobe�   ����  `���  ����*  ����  Qc     �  `���  n���1 1 Qc  ����          -�|  �����  a����  �����  ����  Qb     ��  a����  o���1 1 Qb�  ����          ��  Cor2.   m���r   I���                       �.   a���A   a���0 0                  �.   U���A   U���1 1                   �q   [���c   [���1 1                  2�  y���X  U���                       �  m���'  m���0 0                  �  a���'  a���1 1                   �X  g���J  g���1 1                  ��  Cand2h   �����   ����                       �h   ����v   ����1 1                  �h   ����v   ����0 0                   ��   �����   ����0 0                  ;�f   f����   B���                       �f   Z���t   Z���1 1                  �f   N���t   N���1 1                   ��   T����   T���1 1                  ;�a  �����  ����                       �a  ����o  ����0 0                  �a  ����o  ����0 0                   ��  �����  ����0 0                  ;�e  _����  ;���                       �e  S���s  S���1 1                  �e  G���s  G���1 1                   ��  M����  M���1 1                  -��  ����  n����  ����"  ����  Qa     ��  n����  |���0 0 Qa�  ����          �w  �����  +���                       �w  Q����  Q���0 0                  �w  i����  i���1 1                  ��  �����  ����1 1                  ��  +����  9���1 1                   ��  i����  i���0 0                  ��  Q����  Q���1 1                  -�d   G���x   '���q   Y����   G���  CLK     �n   '���n   5���0 0 CLKb   '���           ��  Cnet1  ��  Csegment�   �����   ����Y��   �����   ����Y��   �����   ����Y��   �����   ���� 	   W�1  Y��   ����   ���Y��   ����   ���Y��   ����   ���Y��   ����   ��� 
   W�1  Y�%  ����%  ����Y�  ����%  ����Y�  ����  ����Y�%  ����%  ����     W�1  Y�%  $���%  ���Y�  ���%  ���Y�  ���  ���Y�%  $���%  $���   $ W�1  Y��  �����  ����Y��  �����  ����Y��  �����  ����Y��  �����  ���� Q  ( W�1  Y�  `���  \���Y�   \���  \���Y��   \����   \���Y�  `���  `���Y��   \���   \���Y�   \���   ����Y�h   ����e   ����Y�e   ����e   ����Y�h   ����h   ����Y��   ����   ����Y�e   �����   ����Y��   $����   ����Y�e  S����  S���Y�e  S���e  S���Y��  S����  $���Y��   $����  $��� / = I   W�1 
 Y��  a����  b���Y�l  b����  b���Y�G  b���G  b���Y��  a����  a���Y�G  b���l  b���Y�l  b���l  u���Y�d   u���l  u���Y�d   u���d   Z���Y�f   Z���d   Z���Y�f   Z���f   Z��� 1 A   W�0  Y��  n����  n���Y��  n����  i���Y��  i����  i���Y��  i����  i���Y��  i����  ����Y�B   �����  ����Y�B   ����B   ����Y�C   ����B   ����Y�h   ����C   ����Y�h   ����h   ����Y��  i����  i���Y��  i����  i��� M >  S W�0  Y��   ����)  ����Y�)  ����)  ����Y��   �����   ����Y�)  ����.   ����Y�.   a���.   ����Y�.   a���.   a��� 4  ? W�1  Y��   T���H  T���Y�H  ����H  T���Y��   T����   T���Y�H  ����   ����Y�   R���   ����Y�   R���.   R���Y�.   U���.   R���Y�.   U���.   U��� 5  C W�1  Y��   \����   [���Y�q   [����   [���Y�q   [���q   [���Y��   \����   \���   6 W�0 
 Y��   D����  D���Y��  f����  D���Y��   D����   D���Y��  f���  f���Y�  b���  f���Y�  b���  b���Y��  f����  f���Y��  f����  ����Y�a  �����  ����Y�a  ����a  ����  E   W�0  Y�G  J���G  ����Y�a  ����G  ����Y�a  ����a  ����Y�G  J���G  J��� F   W�1  Y��  Q����  Q���Y��  Q����  Q���Y��  v����  Q���Y�@  v����  v���Y�W  G���@  G���Y�@  v���@  G���Y�e  G���e  G���Y�e  G���W  G���Y�W  ���W  G���Y�f   N���f   N���Y�f   N���C   N���Y�C   N���C   ���Y�W  ���C   ��� J B  T W�0  Y��  ����A  ����Y�A  ����A  ����Y��  �����  ����Y�A  ����  ����Y�  m���  ����Y�  m���  m��� 8  G W�1  Y��  M���  M���Y�  ����  M���Y��  M����  M���Y�  ����  ����Y�  _���  ����Y�  _���  _���Y�  a���  _���Y�  a���  a��� 9  K W�1  Y�w  i���w  g���Y�X  g���w  g���Y�X  g���X  g���Y�w  i���w  i��� P  : W�0  Y��   D����   (���Y�n   (����   (���Y�L   (���L   (���Y��   D����   D���Y��   (���  (���Y�  J���  (���Y�  J���  J���Y�  (���w  (���Y�w  Q���w  (���Y�w  Q���w  Q���Y�L   (���n   (���Y�n   (���n   '���Y�n   '���n   '���   O V   W�1  Y��  +����  ���Y��  ����  ���Y��  ����  ���Y��  +����  +��� R  , W�Z         17702