2�d d        �  < ��  Cxor2Y  �����  i���                       ��  CpinY  ����l  ����0 0                  �Y  u���l  u���0 0                   ��  {����  {���0 0                  ��  b���   >���                       ��  V����  V���0 0                  ��  J����  J���0 0                   ��  P����  P���0 0                  ��  Cand2�   w���4  S���                       ��   k����   k���0 0                  ��   _����   _���0 0                   �3  e���%  e���0 0                  ��   ���9  ����                       ��   ���  ���0 0                  ��   ����  ����0 0                   �8  ���*  ���0 0                  ��   ����9  ����                       ��   ����  ����0 0                  ��   ����  ����0 0                   �8  ����*  ����0 0                  ��  Cor3(  ���l  ����                       �(  ���;  ���0 0                  �(  
���<  
���0 0                  �(  ����;  ����0 0                   �k  
���]  
���0 0                  ��  Cprobe�  q���  Q����  Q���  ?���  SUM     ��  Q����  _���0 0 SUM�  Q���          �b  +���v  ���_  ����  ����  Cout     �l  ���l  ���0 0 Cout_  ���          ��  Cinput_signalz   �����   x����   �����   ���� X       ��   �����   ����0 0 X�   ����         ��  Csignal    0 &��   0 &��  0 &�X  0 &�   1 &��  1 &��  1 &�x  1 #�w   G����   5����   Y����   G��� Y       ��   >����   >���0 0 Y�   L���         &�    0 &��   0 &��  1 &�X  1 &�   0 &��  0 &��  1 &�x  1 #�w   �����   �����   �����   ���� Cin       ��   �����   ����0 0 Cin�   ����         &�    0 &��   1 &��  0 &�X  1 &�   0 &��  1 &��  1 &�x  0 �� 
 CFullAdder�  �����  6���                       ��  6����  D���Z Z                 ��  6����  D���Z Z                 ��  V����  V���Z Z                   ��  V����  V���X X                  ��  �����  z���X X                  #��  �����  ����                         ��  �����  ����Z Z                   &�    Z #��  ����  ���                         ��  ����  ���Z Z                   &�    Z ��  �����  ����                        ��  �����  ����X X                    ��  v����  V���                        ��  V����  d���X X                    C�  M���r  ����                       �<  ����<  	���0 0                 �P  ����P  	���1 1                 �r  ���d  ���1 1                   �  ���(  ���1 1                  �F  M���F  ?���0 0                  C��  J����  ����                       ��  �����  ���1 1                 ��  �����  ���1 1                 ��  ����  ���1 1                   ��  ����  ���1 1                  ��  J����  <���1 1                  C�%  G���}  ����                       �G  ����G  ���1 1                 �[  ����[  ���1 1                 �}  ���o  ���1 1                   �%  ���3  ���1 1                  �Q  G���Q  9���1 1                  C��  B���	  ����                       ��  �����  ����0 0                 ��  �����  ����1 1                 �	  ����  ���1 1                   ��  ����  ���1 1                  ��  B����  4���0 0                  C�D  ?����  ����                       �f  ����f  ����0 0                 �z  ����z  ����1 1                 ��  ����  ���1 1                   �D  ���R  ���1 1                  �p  ?���p  1���0 0                  C��  ?���"  ����                       ��  �����  ����0 0                 �   ����   ����0 0                 �"  ���  ���1 1                   ��  ����  ���0 0                  ��  ?����  1���1 1                  C�W  >����  ����                       �y  ����y  ����1 1                 ��  �����  ����1 1                 ��  ����  ���0 0                   �W  ���e  ���1 1                  ��  >����  0���0 0                  C�}  �����  1���                       ��  1����  ?���Z Z                 ��  1����  ?���Z Z                 ��  Q����  Q���Z Z                   �}  Q����  Q���X X                  ��  �����  u���X X                  C��  C���>  ����                       �  ����  ����1 1                 �  ����  ����1 1                 �>  ���0  ���1 1                   ��  ����  ���1 1                  �  C���  5���1 1                  C�V  ����  ����                       �x  ����x  ����Z Z                 ��  �����  ����Z Z                 ��  �����  ����Z Z                   �V  ����d  ����X X                  ��  ����   ���X X                  ��  Cswitch�  <����  ����  ����  ���� A7    ��  ����  ���1 0                  ��  ����  ���0                     ��  <����  .���1 0 A7�  ����        ��  =���  ���  ����2  ���� B7    �  ���  ���1                    �  ���  ���0                     �  =���  /���0 0 B7  ����        ��o  <���{  ���e  �����  ���� A6    �o  ���o  ���1                    �{  ���{  ���0                     �u  <���u  .���1 0 A6e  ����        ���  :����  
����  �����  ���� B6    ��  
����  ���1 v                  ��  
����  ���0                     ��  :����  ,���0 0 B6�  ����        ���  ?����  ����  ����  ���� A5    ��  ����  ���1                    ��  ����  ���0                     ��  ?����  1���0 0 A5�  ���        ���  ?���  ����   ���  ���� B5    ��  ����  ���1                    �  ���  ���0                     ��  ?����  1���1 0 B5�   ���        ��_  A���k  ���U  ����v  ���� A4    �_  ���_  ���1                    �k  ���k  ���0                     �e  A���e  3���0 0 A4U  ����        ��x  A����  ���~  �����  ���� B4    �x  ���x  ���1                    ��  ����  ���0                     �~  A���~  3���0 0 B4~  ����        ���  B����  ����  �����  ���� A3    ��  ����   ���1                    ��  ����   ���0                     ��  B����  4���0 0 A3�  ����        ���  A����  ����  ���  ���� B3    ��  ����  ���1                    ��  ����  ���0                     ��  A����  3���0 0 B3�  ���        ��@  D���L  ���5  ���V  ���� A2    �@  ���@  "���1                    �L  ���L  "���0                     �F  D���F  6���1 0 A25  ���        ��Y  D���e  ���\  ���}  ���� B2    �Y  ���Y  "���1                    �e  ���e  "���0                     �_  D���_  6���0 0 B2\  ���        ���  I����  ����  �����  ���� A1    ��  ����  '���1                    ��  ����  '���0                     ��  I����  ;���1 0 A1�  ����        ���  H����  ����  �����  ���� B1    ��  ����  &���1                    ��  ����  &���0                     ��  H����  :���0 0 B1�  ����        ��;  H���G  ���:  ����[  ���� A0    �;  ���;  &���1                    �G  ���G  &���0                     �A  H���A  :���0 0 A0:  ����        ��U  I���a  ���X  ����y  ���� B0    �U  ���U  '���1                    �a  ���a  '���0                     �[  I���[  ;���0 0 B0X  ����        �!  ����e  ~���                       �!  ����4  ����0 0                  �!  ����4  ����1 1                   �d  ����V  ����1 1                  ��  �����  ����                       ��  �����  ����0 0                  ��  �����  ����1 1                   ��  �����  ����1 1                  �  ����L  |���                       �  ����  ����1 1                  �  ����  ����1 1                   �K  ����=  ����0 0                  ��  �����  t���                       ��  �����  ����0 0                  ��  �����  ����1 1                   ��  �����  ����1 1                  ��  ����;  s���                       ��  ����
  ����0 0                  ��  ���
  ���1 1                   �:  ����,  ����1 1                  �l  �����  n���                       �l  ����  ����0 0                  �l  z���  z���1 1                   ��  �����  ����1 1                  ��  ����$  i���                       ��  �����  ����0 0                  ��  u����  u���1 1                   �#  {���  {���1 1                  �`  �����  i���                       �`  ����s  ����0 0                  �`  u���s  u���1 1                   ��  {����  {���1 1                  �  c���  C���                        �  C���  Q���1 1                    �  b����  B���                        ��  B����  P���0 0                    ��  `���  @���                        ��  @����  N���1 1                    �f  `���z  @���                        �p  @���p  N���0 0                    ��  b����  B���                        ��  B����  P���0 0                    �H  g���\  G���                        �R  G���R  U���1 1                    ��  l����  L���                        ��  L����  Z���1 1                    �<  l���P  L���                        �F  L���F  Z���0 0                    ��  0����  ���                        ��  ����  ���1 1                    ���  !���  ����  3���  !��� Cin.    �  ���  ���1                    �  !���  !���0                     ��  ����  ���1 0 Cin.�  3���        : ��  Cnet0  ��  Csegment�   �����   ����	�Y  ����Y  ����	�Y  �����   ����	��   �����   k���	��   k����   k���	��   k����   k���	��   �����   ����	��   �����   ����	��   �����   ����	��   �����   ����	��   �����   ����     % �0  	�Y  u���Y  >���	��   >���Y  >���	�Y  u���Y  u���	��   >����   >���	��   >����   _���	��   _����   _���	��   _����   _���	��   >����   >���	��   >����   ���	��   ����   ���	��   ����   ���	��   ����   ���	��   ����   ���	��   >����   >���     0 �0  	��  V����  V���	��  V����  {���	��  {����  {���	��  {����  {���	��  V����  V���    �0  	�(  ���(  e���	�3  e���(  e���	�3  e���3  e���	�(  ���(  ���    �0  	�(  
���(  ���	�8  ���(  ���	�8  ���8  ���	�(  
���(  
���    �0  	�(  ����(  ����	�8  ����(  ����	�8  ����8  ����	�(  ����(  ����    �0  	��  J����  J���	��  J����  ����	��  �����   ����	��   �����   ����	��   �����   ����	��   �����   ����	��   �����   ����	��   �����   ����	��   �����   ����	��   �����   ����	��   �����   ����	��   �����   ���� 	    : �0  	��  P����  Q���	��  Q����  Q���	��  Q����  Q���	��  P����  P���    
 �0  	�k  
���k  ���	�l  ���k  ���	�l  ���l  ���	�k  
���k  
��� "   �X  	��  �����  ����	��  �����  ����	��  �����  ����	��  �����  ���� Q  I �X  	��  V����  V���	��  V����  V���	��  V����  V��� S  H �Z  	��  6����  ���	��  ����  ���	��  ����  ���	��  6����  6��� E  N �Z  	��  �����  ����	��  �����  ����	��  �����  6���	��  6����  6���	��  6����  6��� F  K �Z  	��  i����  V���	��  V����  V��� G   �1  	��  ����  ���	�  ����  ���	�  ���  ���	��  ����  ��� ]  X �1  	�}  ���}  ���	��  ���}  ���	��  ����  ���	�}  ���}  ��� c  ^ �1  	�	  ���	  ���	�%  ���	  ���	�%  ���%  ���	�	  ���	  ��� i  d �1  	��  ����  ���	��  ����  ���	��  ����  ���	��  ����  ��� o  j �1  	�D  ���"  ���	�D  ���D  ���	�"  ���"  ��� u  p �0  	��  ����  ���	��  ����  ���	��  ����  ���	��  ����  ��� {  v �1  	�>  ���>  ���	�W  ���W  ���	�>  ���>  ���	�>  ���>  ���	�W  ���>  ��� �  | �0  	�  =���  =���	�  ����  =���	�  =���  =���	�  ����!  ����	�!  ����!  ����	�!  ����!  ���� �  � �0  	��  :����  ����	��  :����  :���	��  �����  ����	��  �����  ����	��  �����  ���� �  � �1  	��  ?����  ����	��  ?����  ?���	��  ����  ����	�  ����  ����	�  ����  ���� �  � �0  	�~  A���y  A���	�y  ����y  A���	�~  A���~  A���	�y  �����  ����	��  �����  ����	��  �����  ���� �  � �0  	��  A����  A���	��  �����  A���	��  A����  A���	��  �����  ����	��  �����  ����	��  �����  ���� �  � �0  	�_  D���_  ����	�_  D���_  D���	�_  ����l  ����	�l  ����l  ����	�l  ����l  ���� �  � �0  	��  H����  ����	��  H����  H���	��  �����  ����	��  �����  ����	��  �����  ���� �  � �0  	�[  I���T  I���	�T  ����T  I���	�[  I���[  I���	�T  ����`  ����	�`  ����`  ����	�`  ����`  ���� �  � �Z       �Z       �Z       �1  	�d  ����d  ����	�  ����d  ����	�  ����  ����	�d  ����d  ���� �  � �1  	��  �����  ����	��  �����  ����	��  �����  ����	��  �����  ���� z  � �0  	�K  ����K  ����	�   ����K  ����	�   ����   ����	�K  ����K  ���� t  � �1  	��  �����  ����	�z  �����  ����	�z  ����z  ����	��  �����  ���� n  � �1  	�:  ����:  ����	��  ����:  ����	��  �����  ����	�:  ����:  ���� h  � �1  	��  �����  ����	�[  �����  ����	�[  ����[  ����	��  �����  ���� b  � �1  	�#  {���#  ����	��  ����#  ����	��  �����  ����	�#  {���#  {��� \  � �1  	��  {����  ����	�P  �����  ����	�P  ����P  ����	��  {����  {��� V  � �1  	�  <���  ����	��  <����  <���	�  ����  ����	��  <���  <��� �  � �1  	�u  ����u  <���	�y  ����y  ����	�u  <���u  <���	�y  ����u  ���� y  � �0  	�e  A���e  ����	�f  ����e  ����	�f  ����f  ����	�e  A���e  A��� m  � �0  	��  B����  ����	��  �����  ����	��  �����  ����	��  B����  B��� g  � �1  	�F  D���F  ����	�G  ����F  ����	�G  ����G  ����	�F  D���F  D��� a  � �1  	��  I����  ����	��  �����  ����	��  �����  ����	��  I����  I��� [  � �0  	�A  H���A  ����	�<  ����A  ����	�<  ����<  ����	�A  H���A  H��� U  � �1  	�  C���  C���	�  C���  C��� �  � �0  	��  B����  B���	��  >����  >���	��  B����  B���	��  >����  B��� �  } �1  	��  ?����  @���	��  @����  @���	��  @����  @���	��  ?����  ?��� �  w �0  	�p  @���p  ?���	�p  @���p  @���	�p  ?���p  ?��� �  q �0  	��  B����  B���	��  B����  B��� �  k �1  	�R  G���Q  G���	�R  G���R  G���	�Q  G���Q  G��� �  e �1  	��  J����  L���	��  L����  L���	��  L����  L���	��  J����  J��� �  _ �0  	�F  L���F  M���	�F  L���F  L���	�F  M���F  M���   Y �0  	��  ?����  ����	��  �����  ����	��  �����  ����	��  ?����  ?��� s  � �1  	��  ����  ���	��  ����  ���	��  ����  ���	��  ����  ���  � �1 ! 	�r  ���r  ���	��  ���r  ���	��  ����  V���	�`  V����  V���	��  V���`  V���	�`  V���`  u���	�`  u���`  u���	�p  V����  V���	��  V����  u���	��  u����  u���	��  u����  u���	��  V���p  V���	�p  V���p  z���	�l  z���p  z���	�l  z���l  z���	��  V����  V���	��  V����  ���	��  ����  ���	�  V����  V���	��  V����  ����	��  �����  ����	��  �����  ����	��  V���  V���	�  V���  ����	�  ����  ����	�  V����  V���	��  V����  ����	��  �����  ����	�  V���  ����	�!  ����  ����	�!  ����!  ����	��  ����  ���	��  ����  ���	 W � � � � � � � �    James