2�d d           ��  Cclock'   4���]   "���                
         ��  Cpin]   +���O   +���0 1                  �� 
 CDflipflop�   ����   0���                       ��   V����   V���0 0                  ��   n����   n���1 1                  ��   �����   ����1 1                  ��   0����   >���1 1                   �   n����   n���1 1                  �   V����   V���0 0                  ��  ����C  +���                       ��  Q���  Q���0 0                  ��  i���  i���0 0                  �!  ����!  ����1 1                  �!  +���!  9���1 1                   �C  i���5  i���1 1                  �C  Q���5  Q���0 0                  �S  �����  *���                       �S  P���a  P���0 0                  �S  h���a  h���1 1                  �u  ����u  ����1 1                  �u  *���u  8���1 1                   ��  h����  h���0 0                  ��  P����  P���1 1                  ��  Cswitch�   �����   ����                       ��   �����   ����1                    ��   �����   ����0                     ��   �����   ����1 1                  ��   ����   ���                       ��   ����   ���1                    ��   ����   ���0                     ��   ����   ���1 1                  ��  ����  ����                       ��  �����  ����1                    ��  �����  ����0                     �  �����  ����1 1                  ��  ���  ���                       ��  ����  ���1                    ��  ����  ���0                     �  ���  ���1 1                  �5  ���e  ���                       �5  ���C  ���1                    �5  ���C  ���0                     �e  ���W  ���1 1                  ��  Cor2�   �����   ����                       ��   �����   ����1 1                  ��   �����   ����1 1                   ��   �����   ����1 1                  ��  Cor3h  �����  ����                       �h  ����{  ����0 0                  �h  ����|  ����1 1                  �h  ����{  ����0 0                   ��  �����  ����1 1                  ��  Cand2�  �����  ����                       ��  �����  ����0 0                  ��  �����  ����1 1                   ��  �����  ����0 0                  ;��  ����!  ����                       ��  �����  ����0 0                  ��  �����  ����1 1                   �!  ����  ����0 0                  ;��  ����!  c���                       ��  {����  {���1 1                  ��  o����  o���1 1                   �!  u���  u���1 1                  ��  Cand3�  :���  ���                       ��  4����  4���1 1                  ��  (����  (���0 0                  ��  ����  ���0 0                   �  (���  (���0 0                  ��  Cprobe  ����,  q���%  ����G  ����  Qc     �"  q���"  ���1 1 Qc%  ����          N�e  ����y  i���r  �����  ����  Qb     �o  i���o  w���1 1 Qbr  ����          N��  �����  g����  �����  ����  Qa     ��  g����  u���0 0 Qa�  ����          �+  ����[  ����                       �+  ����9  ����1                    �+  ����9  ����0                     �[  ����M  ����1 1                  �e  �����  ����                       �e  ����s  ����1                    �e  ����s  ����0                     ��  �����  ����1 1                   ��  Cnet1  ��  Csegment�   0����   ���_��   ����   ���_��   ����   ���_��   0����   0��� 
  # ]�1  _��   �����   ����_��   �����   ����_��   �����   ����_��   �����   ���� 	   ]�1  _�"  q���"  n���_�  n���"  n���_�   n���   n���_�"  q���"  q���_�   n���  n���_�  n���  4���_��  4���  4���_��  4����  4��� P J   ]�1  _�g  i���o  i���_�C  i���C  i���_�o  i���o  i���_�C  i���\  i���_�\  i���\  ����_��   �����   ����_��   �����   ����_��   �����   ����_��   ����\  ����_�\  i���g  i���_�g  i���g  {���_��  {���g  {���_��  {����  {��� R 2 E   ]�1  _�!  ����!  ����_�  ����!  ����_�  ����  ����_�!  ����!  ����   ' ]�1  _�!  +���!  ���_�  ���!  ���_�  ���  ���_�!  +���!  +���   + ]�1  _�u  ����u  ����_�[  ����u  ����_�u  ����u  ����_�[  ����[  ����   X ]�1  _�u  *���u  ���_�e  ���u  ���_�e  ���e  ���_�u  *���u  *���   / ]�0  _��  g����  g���_��  g����  h���_��  h����  h���_��  h����  h���_��  h����  h���_��  h����  h���_��  �����  h���_��  ����  ���_��  ����  ���_��  �����  ���_��  �����  ����_��  �����  ���� T L   ]�1  _��   ����K  ����_�K  ����K  ����_��   �����   ����_�K  �����   ����_��   n����   ����_��   n����   n���   4 ]�0 
 _��   V����   +���_�]   +����   +���_�]   +���]   +���_��   V����   V���_��   +����  +���_��  Q����  +���_��  Q����  Q���_��  +���S  +���_�S  P���S  +���_�S  P���S  P���      ]�0  _��  �����  ����_��  �����  ����_��  �����  ����_��  �����  ����_��  i����  ����_��  i����  i���   ? ]�0 
 _��  �����  ����_��  �����  ����_��  �����  ����_�$  ����C  ����_�C  Q���C  ����_�C  Q���C  Q���_��  ����$  ����_�$  ����$  (���_��  (���$  (���_��  (����  (��� = K   ]�1  _��  �����  ����_��  �����  ����_��  �����  ����_�,  �����  ����_��  P����  ����_��  P����  P���_��  �����  ����_��  �����  ����_��  �����  ����_��  �����  ����_��  �����  o���_��  o����  o���_��  o����  o���_��  ����,  ����_�,  ����,  E���_��   �����   ����_��   �����   ����_��   E����   ����_��   E���,  E��� > B F 3   ]�0  _�   V���   ����_��  ����   ����_��  �����  ����_�   V���   V��� A   ]�0  _�h  ����h  ����_�!  ����h  ����_�!  ����!  ����_�h  ����h  ���� 7  C ]�1  _�!  u���!  ����_�h  ����!  ����_�h  ����h  ����_�!  u���!  u��� 8  G ]�0  _�h  ����1  ����_�1  (���1  ����_�h  ����h  ����_�1  (���  (���_�  (���  (��� 9  M ]�1  _��  �����  ����_��  �����  ����_��  �����  ����_��  ����S  ����_�S  h���S  ����_�S  h���S  h���   :   17702